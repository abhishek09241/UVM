module hello;
	initial
		$display("Hello , Welecom to My Git Hub in Learning UVM",);

endmodule : hello